LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY Forwarding IS
PORT (
EXMEMRegWrite, MEMWBRegWrite : IN STD_LOGIC;
EXMEMRD, IDEXRS, IDEXRT, MEMWBRD : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
fwdA, fwdB : OUT STD_LOGIC_VECTOR(1 DOWNTO 0));
END Forwarding;

ARCHITECTURE structural OF Forwarding IS
SIGNAL notZero, eqRS_EXMEM,eqRT_EXMEM, eqRS_MEMWB, eqRT_MEMWB : STD_LOGIC;

BEGIN
    eqRS_EXMEM <= (EXMEMRD(4) XNOR IDEXRS(4)) AND (EXMEMRD(3) XNOR IDEXRS(3)) AND (EXMEMRD(2) XNOR IDEXRS(2)) AND (EXMEMRD(1) XNOR IDEXRS(1)) AND (EXMEMRD(0) XNOR IDEXRS(0));
    eqRT_EXMEM <= (EXMEMRD(4) XNOR IDEXRT(4)) AND (EXMEMRD(3) XNOR IDEXRT(3)) AND (EXMEMRD(2) XNOR IDEXRT(2)) AND (EXMEMRD(1) XNOR IDEXRT(1)) AND (EXMEMRD(0) XNOR IDEXRT(0));
    eqRS_MEMWB <= (MEMWBRD(4) XNOR IDEXRS(4)) AND (MEMWBRD(3) XNOR IDEXRS(3)) AND (MEMWBRD(2) XNOR IDEXRS(2)) AND (MEMWBRD(1) XNOR IDEXRS(1)) AND (MEMWBRD(0) XNOR IDEXRS(0));
    eqRT_MEMWB <= (MEMWBRD(4) XNOR IDEXRT(4)) AND (MEMWBRD(3) XNOR IDEXRT(3)) AND (MEMWBRD(2) XNOR IDEXRT(2)) AND (MEMWBRD(1) XNOR IDEXRT(1)) AND (MEMWBRD(0) XNOR IDEXRT(0));
	 notZero <= EXMEMRegWrite AND (EXMEMRD(4)Or EXMEMRD(3)Or EXMEMRD(2)Or EXMEMRD(1)Or EXMEMRD(0));
	 
    fwdA(1)<= notZero AND eqRS_EXMEM;
	 fwdA(0)<= notZero AND eqRS_MEMWB;
    fwdB(1)<= notZero AND eqRT_EXMEM;
	 fwdB(0)<= notZero AND eqRT_MEMWB;
	 
END structural;